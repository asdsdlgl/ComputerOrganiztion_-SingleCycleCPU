// Controller

module Controller ( opcode,
					funct,
					ALUOp,
					RegWrite,
					Branch,
					Jr,
					Jump,
					Jal,
					MemWrite,
					MemToReg,
					RegDst,
					Signextend
					);

	input  [5:0] opcode;
	input  [5:0] funct;
	output [3:0] ALUOp;
	output RegWrite;
	output MemWrite;
	output MemToReg;
	output Branch;
	output Jr;
	output Jump;
	output Jal;
	output RegDst;
	output Signextend;
	reg [3:0] ALUOp;
	reg RegWrite;
	reg MemToReg;
	reg MemWrite;
	reg Branch;
	reg Jr;
	reg Jump;
	reg Jal;
	reg RegDst;
	reg Signextend;
	always @(*)	
		begin
		RegWrite = 0;
		MemToReg = 0;
		MemWrite = 0;
		Branch = 0;
		Jr = 0;
		Jump = 0;
		Jal = 0;
		RegDst = 0;
		Signextend = 0;
		case(opcode)
			6'b000000:
				begin
				case(funct)
					6'b100000:
					begin
						ALUOp = 4'b0000;//add
						RegWrite = 1;
					end
					6'b100010:
					begin
						ALUOp = 4'b0001;//sub
						RegWrite = 1;
					end
					6'b100100:
					begin
						ALUOp= 4'b0010;//and
						RegWrite = 1;
					end
					6'b100101:
					begin
						ALUOp = 4'b0011;//or
						RegWrite = 1;
					end
					6'b100110:
					begin
						ALUOp = 4'b0100;//xor
						RegWrite = 1;
					end
					6'b100111:
					begin
						ALUOp = 4'b0101;//nor
						RegWrite = 1;
					end
					6'b101010:
					begin
						ALUOp = 4'b0110;//less
						RegWrite = 1;
					end
					6'b000000:
					begin
						ALUOp = 4'b0111;//left shift
						RegWrite = 1;
					end
					6'b000010:
					begin
						ALUOp = 4'b1000;//right shift
						RegWrite = 1;
					end
					6'b001000://JR
					begin
						Jr = 1;
					end
					6'B001001://Jalr
					begin
						Jal = 1;
						Jr = 1;
					end
					//6'b001000:ALUOp = 4'b1001;//beq
					//6'b100000:ALUOp = 4'b1010;//bne
				endcase
				end
			6'b001000:
			begin
				ALUOp = 4'b0000;//addi
				RegWrite = 1;
				RegDst = 1;
			end
			6'b001100:
			begin
				ALUOp = 4'b0010;//andi
				RegWrite = 1;
				RegDst = 1;
			end
			6'b001010:
			begin
				ALUOp = 4'b0110;//slti
				RegWrite = 1;
				RegDst = 1;
			end
			6'b001101:
			begin
				ALUOp = 4'b0011;//ori
				RegWrite = 1;
				RegDst = 1;
			end
			6'b000100:
			begin
				ALUOp = 4'b1001;//equal
				Branch = 1;
			end
			6'b000101:
			begin
				ALUOp = 4'b1010;//bne
				Branch = 1;
			end
			6'b100011:
			begin
				ALUOp = 4'b0000;//lw->add
				RegWrite = 1;
				MemToReg = 1;
				RegDst = 1;
			end
			6'b101011:
			begin
				ALUOp = 4'b0000;//sw->add
				MemWrite = 1;
				RegDst = 1;
			end
			6'b100001:
			begin
				ALUOp = 4'b0000;//lh->add
				Signextend = 1;
				RegWrite = 1;
				MemToReg = 1;
				RegDst = 1;
			end
			6'b101001:
			begin
				ALUOp = 4'b0000;//sh->add
				Signextend = 1;
				MemWrite = 1;
				RegDst = 1;
			end
			6'b000010://jump
			begin
				Jump = 1;
			end
			6'b000011://jal
			begin
				Jump = 1;
				Jal = 1;
				RegWrite = 1;
			end
		endcase
		end
	
endmodule




